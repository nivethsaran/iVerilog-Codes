module months_tb;
reg i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11;
wire o0,o1,o2;
months m1(i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,o0,o1,o2);
initial
begin
    $monitor("%b  %b  %b  %b  %b  %b  %b  %b  %b  %b  %b   %b   %b  %b  %b ",i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,o0,o1,o2);
    $display("i0 i1 i2 i3 i4 i5 i6 i7 i8 i9 i10 i11 o0 o1 o2");
i0=1'b1;
i1=1'b0;
i2=1'b0;
i3=1'b0;
i4=1'b0;
i5=1'b0;
i6=1'b0;
i7=1'b0;
i8=1'b0;
i9=1'b0;
i10=1'b0;
i11=1'b0;
#5
i0=1'b0;
i1=1'b1;
i2=1'b0;
i3=1'b0;
i4=1'b0;
i5=1'b0;
i6=1'b0;
i7=1'b0;
i8=1'b0;
i9=1'b0;
i10=1'b0;
i11=1'b0;
#5
i0=1'b0;
i1=1'b0;
i2=1'b1;
i3=1'b0;
i4=1'b0;
i5=1'b0;
i6=1'b0;
i7=1'b0;
i8=1'b0;
i9=1'b0;
i10=1'b0;
i11=1'b0;
#5
i0=1'b0;
i1=1'b0;
i2=1'b0;
i3=1'b1;
i4=1'b0;
i5=1'b0;
i6=1'b0;
i7=1'b0;
i8=1'b0;
i9=1'b0;
i10=1'b0;
i11=1'b0;
#5
i0=1'b0;
i1=1'b0;
i2=1'b0;
i3=1'b0;
i4=1'b1;
i5=1'b0;
i6=1'b0;
i7=1'b0;
i8=1'b0;
i9=1'b0;
i10=1'b0;
i11=1'b0;
#5
i0=1'b0;
i1=1'b0;
i2=1'b0;
i3=1'b0;
i4=1'b0;
i5=1'b1;
i6=1'b0;
i7=1'b0;
i8=1'b0;
i9=1'b0;
i10=1'b0;
i11=1'b0;
#5
i0=1'b0;
i1=1'b0;
i2=1'b0;
i3=1'b0;
i4=1'b0;
i5=1'b0;
i6=1'b1;
i7=1'b0;
i8=1'b0;
i9=1'b0;
i10=1'b0;
i11=1'b0;
#5
i0=1'b0;
i1=1'b0;
i2=1'b0;
i3=1'b0;
i4=1'b0;
i5=1'b0;
i6=1'b0;
i7=1'b1;
i8=1'b0;
i9=1'b0;
i10=1'b0;
i11=1'b0;
#5
i0=1'b0;
i1=1'b0;
i2=1'b0;
i3=1'b0;
i4=1'b0;
i5=1'b0;
i6=1'b0;
i7=1'b0;
i8=1'b1;
i9=1'b0;
i10=1'b0;
i11=1'b0;
#5
i0=1'b0;
i1=1'b0;
i2=1'b0;
i3=1'b0;
i4=1'b0;
i5=1'b0;
i6=1'b0;
i7=1'b0;
i8=1'b0;
i9=1'b1;
i10=1'b0;
i11=1'b0;
#5
i0=1'b0;
i1=1'b0;
i2=1'b0;
i3=1'b0;
i4=1'b0;
i5=1'b0;
i6=1'b0;
i7=1'b0;
i8=1'b0;
i9=1'b0;
i10=1'b1;
i11=1'b0;
#5
i0=1'b0;
i1=1'b0;
i2=1'b0;
i3=1'b0;
i4=1'b0;
i5=1'b0;
i6=1'b0;
i7=1'b0;
i8=1'b0;
i9=1'b0;
i10=1'b0;
i11=1'b1;
end
endmodule
