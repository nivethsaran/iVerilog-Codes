module hexto7seg_tb;

    reg [15:0] hex;
    wire [6:0] seg;

hexto7seg hexto7seg1(.hex(hex),.seg(seg));

initial 
begin
$monitor("%b %b",hex,seg);
        
hex=16'b1000000000000000;
#10
hex=16'b0100000000000000;
#10
hex=16'b0010000000000000;
#10
hex=16'b0001000000000000;
#10
hex=16'b0000100000000000;
#10
hex=16'b0000010000000000;
#10
hex=16'b0000001000000000;
#10
hex=16'b0000000100000000;
#10
hex=16'b0000000010000000;
#10
hex=16'b0000000001000000;
#10
hex=16'b0000000000100000;
#10
hex=16'b0000000000010000;
#10
hex=16'b0000000000001000;
#10
hex=16'b0000000000000100;
#10
hex=16'b0000000000000010;
#10
hex=16'b0000000000000001;

end
      
endmodule