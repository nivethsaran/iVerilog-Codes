module hexto7seg(hex,seg);
input  [15:0]hex;
output [6:0]seg;
reg [6:0]seg;
always @(hex)
begin
case (hex)
16'b1000000000000000 : seg = 7'b1111110;
16'b0100000000000000 : seg = 7'b0110000; 
16'b0010000000000000 : seg = 7'b1101101;
16'b0001000000000000 : seg = 7'b1111001;
16'b0000100000000000 : seg = 7'b0110011;
16'b0000010000000000 : seg = 7'b1011011;
16'b0000001000000000 : seg = 7'b1011111;
16'b0000000100000000 : seg = 7'b1110000;
16'b0000000010000000 : seg = 7'b1111111;
16'b0000000001000000 : seg = 7'b1111011;
16'b0000000000100000 : seg = 7'b1110111; 
16'b0000000000010000 : seg = 7'b0011111;
16'b0000000000001000 : seg = 7'b1001110;
16'b0000000000000100 : seg = 7'b0111101;
16'b0000000000000010 : seg = 7'b1001111;
16'b0000000000000001 : seg = 7'b1000111;
endcase
 end
endmodule
